library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.P65816_pkg.all;

entity MCode is
    port( 
        CLK		: in std_logic;
		  RST_N	: in std_logic;
		  EN		: in std_logic;
        IR		: in std_logic_vector(7 downto 0);
        STATE	: in unsigned(3 downto 0);
        M		: out MCode_r
    );
end MCode;

architecture rtl of MCode is

	type MicroInst_t is array(0 to 2047) of MicroInst_r;
	constant  M_TAB: MicroInst_t := (
	-- 00 BRK
	("111","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['PC++'] 
	("000","010","00","000","00","00","00000000","000","011","000","00","000000","00000","01","110","10"),-- ['PBR->[00:SP--]']
	("000","010","00","000","00","00","00000000","000","011","000","00","000000","00000","10","010","10"),-- ['PCH->[00:SP--]'] 
	("000","010","00","000","00","00","00000000","000","011","000","00","000000","00000","01","010","10"),-- ['PCL->[00:SP--]'] 
	("000","010","00","010","00","00","00000000","000","011","000","00","000000","00000","01","100","10"),-- ['P->[00:SP--]']
	("000","100","00","000","00","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:VECT+0]->DR']
	("010","100","01","000","00","00","00000000","010","000","000","10","000000","00000","10","000","10"),-- ['[00:VECT+1]:DR->PC', '00->PBR', '1->I']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 01 ORA (DP,X)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[DX+1]->AAH']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00100","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']  
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00100","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 02 COP
	("111","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['PC++'] 
	("000","010","00","000","00","00","00000000","000","011","000","00","000000","00000","01","110","10"),-- ['PBR->[00:SP--]']
	("000","010","00","000","00","00","00000000","000","011","000","00","000000","00000","10","010","10"),-- ['PCH->[00:SP--]'] 
	("000","010","00","000","00","00","00000000","000","011","000","00","000000","00000","01","010","10"),-- ['PCL->[00:SP--]'] 
	("000","010","00","010","00","00","00000000","000","011","000","00","000000","00000","01","100","10"),-- ['P->[00:SP--]']
	("000","100","00","000","00","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:VECT+0]->DR']
	("010","100","01","000","00","00","00000000","010","000","000","10","000000","00000","10","000","10"),-- ['[00:VECT+1]:DR->PC', '00->PBR', '1->I']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 03 ORA S
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['SPH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00100","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']   
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00100","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 04 TSB DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("110","011","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:DX+0]->TL'] 
	("000","011","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[00:DX+1]->TH'] 
	("110","011","01","001","10","00","00000000","000","000","000","00","000100","01111","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","011","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[00:DX+1]']
	("010","011","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[00:DX+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 05 ORA DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00100","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']   
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00100","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 06 ASL DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("110","011","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:DX+0]->TL'] 
	("000","011","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[00:DX+1]->TH'] 
	("110","011","01","001","10","00","00000000","000","000","000","00","000100","01010","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","011","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[00:DX+1]']
	("010","011","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[00:DX+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 07 ORA [DP]
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("000","011","10","000","00","00","00000001","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00100","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00100","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 08 PHP
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("010","010","00","000","00","00","00000000","000","011","000","00","000000","00000","01","100","10"),-- ['P->[00:SP--]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 09 ORA IMM
	("100","000","00","001","00","00","00000000","001","000","101","00","000000","00100","01","000","01"),-- ['ALU([PBR:PC])->AL', '[PBR:PC]->DR', 'PC++', 'Flags'] 
	("010","000","00","001","00","00","00000000","001","000","101","00","000001","00100","10","000","01"),-- ['ALU([PBR:PC]:DR)->A', 'PC++', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 0A ASL A
	("010","000","00","001","00","00","00000000","000","000","101","00","000010","01010","11","000","00"),-- ['ALU(A)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 0B PHD
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("000","010","00","000","00","00","00000000","000","011","000","00","011000","00000","10","101","10"),-- ['DH->[00:SP]', 'SP--']
	("010","010","00","000","00","00","00000000","000","011","000","00","011000","00000","01","101","10"),-- ['DL->[00:SP]', 'SP--']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 0C TSB ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++'] 
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++'] 
	("110","001","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[DBR:AA+0]->TL'] 
	("000","001","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[DBR:AA+1]->TH'] 
	("110","001","01","001","10","00","00000000","000","000","000","00","000100","01111","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","001","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[DBR:AA+1]']
	("010","001","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[DBR:AA+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 0D ORA ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00100","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags'] 
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00100","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 0E ASL ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++'] 
	("110","001","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[DBR:AA+0]->TL'] 
	("000","001","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[DBR:AA+1]->TH'] 
	("110","001","01","001","10","00","00000000","000","000","000","00","000100","01010","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","001","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[DBR:AA+1]']
	("010","001","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[DBR:AA+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 0F ORA LONG
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("000","000","00","000","00","00","00000001","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'PC++']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00100","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags'] 
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00100","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 10 BPL
	("010","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->DR', 'PC++'] 
	("011","000","00","000","00","00","00000000","100","000","000","00","000000","00000","00","000","00"),-- ['PC+DR->PC']
	("010","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- [] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 11 ORA (DP),Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB']
	("001","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH','AAL+YL->AAL']
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00100","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00100","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 12 ORA (DP)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00100","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']  
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00100","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 13 ORA (S),Y
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['SPH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB']
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL']
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00100","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00100","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 14 TRB DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("110","011","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:DX+0]->TL'] 
	("000","011","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[00:DX+1]->TH'] 
	("110","011","01","001","10","00","00000000","000","000","000","00","000100","01110","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","011","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[00:DX+1]']
	("010","011","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[00:DX+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 15 ORA DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+Carry->DX'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00100","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00100","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 16 ASL DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("110","011","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:DX+0]->TL'] 
	("000","011","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[00:DX+1]->TH'] 
	("110","011","01","001","10","00","00000000","000","000","000","00","000100","01010","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","011","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[00:DX+1]']
	("010","011","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[00:DX+0]']
	-- 17 ORA [DP],Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH','AAL+YL->AAL']
	("000","011","10","000","00","01","00000101","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB','AAH+YH+AALCarry->AAH']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00100","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00100","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 18 CLC
	("010","000","00","100","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- ['Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 19 ORA ABS,Y
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'DBR->AB', 'PC++']
	("001","000","00","000","00","01","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++'] 
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00100","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags'] 
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00100","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 1A INC A
	("010","000","00","001","00","00","00000000","000","000","101","00","000010","00011","11","000","00"),-- ['ALU(A)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 1B TCS
	("010","000","00","000","00","00","00000000","000","100","000","00","000000","00000","00","000","00"),-- ['A->S'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 1C TRB ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++'] 
	("110","001","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[DBR:AA+0]->TL'] 
	("000","001","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[DBR:AA+1]->TH'] 
	("110","001","01","001","10","00","00000000","000","000","000","00","000100","01110","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","001","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[DBR:AA+1]']
	("010","001","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[DBR:AA+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 1D ORA ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'DBR->AB', 'PC++']
	("001","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH']  
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00100","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags'] 
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00100","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 1E ASL ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'DBR->AB', 'PC++']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("110","101","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[AB:AA+0]->TL'] 
	("000","101","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[AB:AA+1]->TH'] 
	("110","101","01","001","10","00","00000000","000","000","000","00","000100","01010","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","101","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[AB:AA+1]']
	("010","101","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[AB:AA+0]']
	-- 1F ORA LONG,X
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++'] 
	("000","000","00","000","00","00","00000101","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'AAH+XH/YH+AALCarry->AAH', 'PC++']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00100","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags'] 
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00100","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 20 JSR ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL, 'PC++'] 
	("000","000","00","000","00","00","00001000","000","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH'] 
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("000","010","00","000","00","00","00000000","000","011","000","00","000000","00000","10","010","10"),-- ['PCH->[00:SP]', 'SP--'] 
	("010","010","00","000","00","00","00000000","110","011","000","00","000000","00000","01","010","10"),-- ['PCL->[00:SP]', 'SP--', 'AA->PC'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 21 AND (DP,X)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00101","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']  
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00101","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 22 JSR LONG
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++'] 
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++'] 
	("000","010","00","000","00","00","00000000","000","011","000","00","000000","00000","00","110","10"),-- ['PBR->[00:SP]', 'SP--'] 
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("000","000","00","000","00","00","00000000","000","000","000","10","000000","00000","00","000","01"),-- ['[PBR:PC]->PBR'] 
	("000","010","00","000","00","00","00000000","000","011","000","00","000000","00000","10","010","10"),-- ['PCH->[00:SP]', 'SP--'] 
	("010","010","00","000","00","00","00000000","110","011","000","00","000000","00000","01","010","10"),-- ['PCL->[00:SP]', 'SP--', 'AA->PC'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 23 AND S
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['SPH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00101","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']   
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00101","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 24 BIT DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","001","00","000000","01001","01","000","10"),-- ['ALU([00:DX+0])', '[00:DX+0]->DR', 'Flags']   
	("010","011","01","001","00","00","00000000","000","000","001","00","000001","01001","10","000","10"),-- ['ALU([00:DX+1]:DR)', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 25 AND DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00101","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']   
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00101","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 26 ROL DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("110","011","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:DX+0]->TL'] 
	("000","011","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[00:DX+1]->TH'] 
	("110","011","01","001","10","00","00000000","000","000","000","00","000100","01100","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","011","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[00:DX+1]']
	("010","011","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[00:DX+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 27 AND [DP]
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("000","011","10","000","00","00","00000001","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00101","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00101","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 28 PLP
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("000","000","00","000","00","00","00000000","000","001","000","00","000000","00000","00","000","00"),-- ['SP++']
	("010","010","00","011","00","00","00000000","000","000","000","00","000000","00000","00","000","10"),-- ['[SP]->P', 'Flags']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 29 AND IMM
	("100","000","00","001","00","00","00000000","001","000","101","00","000000","00101","01","000","01"),-- ['ALU([PBR:PC])->AL', '[PBR:PC]->DR', 'PC++', 'Flags'] 
	("010","000","00","001","00","00","00000000","001","000","101","00","000001","00101","10","000","01"),-- ['ALU([PBR:PC]:DR)->A', 'PC++', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 2A ROL A
	("010","000","00","001","00","00","00000000","000","000","101","00","000010","01100","11","000","00"),-- ['ALU(A)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 2B PLD
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("000","000","00","000","00","00","00000000","000","001","000","00","000000","00000","00","000","00"),-- ['SP++']
	("000","010","00","000","00","00","00000000","000","001","000","00","000000","00000","01","000","10"),-- ['[00:SP++]->DR']
	("010","010","00","001","00","00","00000000","000","000","000","01","000001","00001","10","000","10"),-- ['ALU([00:SP]:DR)->D', 'Flags']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 2C BIT ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","001","00","00","00000000","000","000","001","00","000000","01001","01","000","10"),-- ['ALU([DBR:AA+0])', '[DBR:AA+0]->DR'] 
	("010","001","01","001","00","00","00000000","000","000","001","00","000001","01001","10","000","10"),-- ['ALU([DBR:AA+1]:DR)'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 2D AND ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00101","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR'] 
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00101","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 2E ROL ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++'] 
	("110","001","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[DBR:AA+0]->TL'] 
	("000","001","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[DBR:AA+1]->TH'] 
	("110","001","01","001","10","00","00000000","000","000","000","00","000100","01100","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","001","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[DBR:AA+1]']
	("010","001","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[DBR:AA+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 2F AND LONG
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("000","000","00","000","00","00","00000001","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'PC++']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00101","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags'] 
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00101","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A, 'Flags''] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 30 BMI
	("010","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->DR', 'PC++'] 
	("011","000","00","000","00","00","00000000","100","000","000","00","000000","00000","00","000","00"),-- ['PC+DR->PC']
	("010","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- [] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 31 AND (DP),Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB']
	("001","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL ']
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00101","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00101","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 32 AND (DP)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00101","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']  
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00101","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 33 AND (S),Y
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DX', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB'] 
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+Y->AAL'] 
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00101","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00101","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 34 BIT DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+Carry->DX'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("100","011","00","001","00","00","00000000","000","000","001","00","000000","01001","01","000","10"),-- ['ALU([00:DX+0]', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","001","00","000001","01001","10","000","10"),-- ['ALU([00:DX+1]', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 35 AND DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+Carry->DX'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00101","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']   
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00101","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 36 ROL DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("110","011","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:DX+0]->TL'] 
	("000","011","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[00:DX+1]->TH'] 
	("110","011","01","001","10","00","00000000","000","000","000","00","000100","01100","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","011","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[00:DX+1]']
	("010","011","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[00:DX+0]']
	-- 37 AND [DP],Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH,AAL+Y->AAL']
	("000","011","10","000","00","01","00000101","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB','AAH+YH+AALCarry->AAH']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00101","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00101","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 38 SEC
	("010","000","00","100","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- ['Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 39 AND ABS,Y
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'DBR->AB', 'PC++']
	("001","000","00","000","00","01","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++'] 
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00101","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00101","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 3A DEC A
	("010","000","00","001","00","00","00000000","000","000","101","00","000010","00010","11","000","00"),-- ['ALU(A)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 3B TSC
	("010","000","00","001","00","00","00000000","000","000","101","00","101010","00001","11","000","00"),-- ['ALU(SP)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 3C BIT ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("001","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","001","00","000000","01001","01","000","10"),-- ['ALU([AB:AA+0])', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","001","00","000001","01001","10","000","10"),-- ['ALU([AB:AA+1])' 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 3D AND ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'DBR->AB', 'PC++']
	("001","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00101","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00101","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']   
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 3E ROL ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'DBR->AB', 'PC++']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH''] 
	("110","101","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[AB:AA+0]->TL'] 
	("000","101","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[AB:AA+1]->TH'] 
	("110","101","01","001","10","00","00000000","000","000","000","00","000100","01100","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","101","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[AB:AA+1]']
	("010","101","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[AB:AA+0]']
	-- 3F AND LONG,X
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL', 'PC++'] 
	("000","000","00","000","00","00","00000101","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'AAH+XH/YH+AALCarry->AAH', 'PC++']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00101","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00101","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 40 RTI
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("000","000","00","000","00","00","00000000","000","001","000","00","000000","00000","00","000","00"),-- ['SP++']
	("000","010","00","011","00","00","00000000","000","001","000","00","000000","00000","00","000","10"),-- ['[00:SP]->P', 'SP++']
	("000","010","00","000","00","00","00000000","000","001","000","00","000000","00000","00","000","10"),-- ['[00:SP]->DR', 'SP++']
	("111","010","00","000","00","00","00000000","010","001","000","00","000000","00000","00","000","10"),-- ['[00:SP]:DR->PC', 'SP++']
	("010","010","00","000","00","00","00000000","000","000","000","10","000000","00000","00","000","10"),-- ['[00:SP]->PBR']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 41 EOR (DP,X)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00110","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']  
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00110","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 42 WDM
	("010","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['PC++'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 43 EOR S
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00110","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']   
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00110","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 44 MVP
	("000","000","00","000","00","00","00000000","001","000","000","11","000000","00000","00","000","01"),-- ['[PBR:PC]->DBR', 'PC++'] 
	("000","000","00","000","00","10","00000001","001","000","110","00","001010","00010","11","000","01"),-- ['[PBR:PC]->ABR', 'PC++', 'X->AA', 'X-1->X'] 
	("000","101","00","000","00","11","00000000","000","000","111","00","010010","00010","11","000","10"),-- ['[ABR:AA]->DR', 'Y->AA', 'Y-1->Y'] 
	("000","001","00","000","00","00","00000000","000","000","000","00","000000","00000","10","110","10"),-- ['DR->[DBR:AA]'] 
	("000","001","00","000","00","00","00000000","111","000","101","00","000101","10000","11","000","00"),-- ['ALU(A)->A', 'PC-3->PC'] 
	("010","001","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- [] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 45 EOR DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00110","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']   
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00110","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 46 LSR DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("110","011","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:DX+0]->TL'] 
	("000","011","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[00:DX+1]->TH'] 
	("110","011","01","001","10","00","00000000","000","000","000","00","000100","01011","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","011","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[00:DX+1]']
	("010","011","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[00:DX+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 47 EOR [DP]
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("000","011","10","000","00","00","00000001","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00110","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']   
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00110","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 48 PHA
	("110","000","00","000","00","00","00000000","000","000","001","00","000000","00000","00","000","00"),-- []
	("000","010","00","000","00","00","00000000","000","011","001","00","000000","00000","10","101","10"),-- ['AH->[00:SP]', 'SP--']
	("010","010","00","000","00","00","00000000","000","011","001","00","000000","00000","01","101","10"),-- ['AL->[00:SP]', 'SP--']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 49 EOR IMM
	("100","000","00","001","00","00","00000000","001","000","101","00","000000","00110","01","000","01"),-- ['ALU([PBR:PC])->AL', '[PBR:PC]->DR', 'PC++', 'Flags'] 
	("010","000","00","001","00","00","00000000","001","000","101","00","000001","00110","10","000","01"),-- ['ALU([PBR:PC]:DR)->A', 'PC++', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 4A LSR A
	("010","000","00","001","00","00","00000000","000","000","101","00","000010","01011","11","000","00"),-- ['ALU(REG+1)->REG', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 4B PHK
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("010","010","00","000","00","00","00000000","000","011","000","00","110000","00000","01","101","10"),-- ['PBR->[00:SP]', 'SP--']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 4C JMP ABS
	("000","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->DR', 'PC++'] 
	("010","000","00","000","00","00","00000000","010","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]:DR->PC'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 4D EOR ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++'] 
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00110","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags'] 
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00110","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 4E LSR ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++'] 
	("110","001","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[DBR:AA+0]->TL'] 
	("000","001","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[DBR:AA+1]->TH'] 
	("110","001","01","001","10","00","00000000","000","000","000","00","000100","01011","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","001","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[DBR:AA+1]']
	("010","001","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[DBR:AA+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 4F EOR LONG
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++'] 
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("000","000","00","000","00","00","00000001","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'PC++']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00110","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00110","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 50 BVC
	("010","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->DL', 'PC++'] 
	("011","000","00","000","00","00","00000000","100","000","000","00","000000","00000","00","000","00"),-- ['PC+DL->PC']
	("010","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- ['NOP'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 51 EOR (DP),Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB']
	("001","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL ']
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00110","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00110","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 52 EOR (DP)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- [00:DX+0]->AAL
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- [00:DX+1]->AAH
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00110","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']  
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00110","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 53 EOR (S),Y
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB']
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL ']
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00110","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']   
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00110","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 54 MVN
	("000","000","00","000","00","00","00000000","001","000","000","11","000000","00000","00","000","01"),-- ['[PBR:PC]->DBR', 'PC++'] 
	("000","000","00","000","00","10","00000001","001","000","110","00","001010","00011","11","000","01"),-- ['[PBR:PC]->ABR', 'PC++', 'X->AA', 'X+1->X'] 
	("000","101","00","000","00","11","00000000","000","000","111","00","010010","00011","11","000","10"),-- ['[ABR:AA]->DR', 'Y->AA', 'Y+1->Y'] 
	("000","001","00","000","00","00","00000000","000","000","000","00","000000","00000","10","110","10"),-- ['DR->[DBR:AA]'] 
	("000","001","00","000","00","00","00000000","111","000","101","00","000101","10000","11","000","00"),-- ['ALU(A-1)->A','PC-3->PC'] 
	("010","001","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- [] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 55 EOR DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+Carry->DX'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00110","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags'] 
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00110","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 56 LSR DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("110","011","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:DX+0]->TL'] 
	("000","011","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[00:DX+1]->TH'] 
	("110","011","01","001","10","00","00000000","000","000","000","00","000100","01011","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","011","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[00:DX+1]']
	("010","011","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[00:DX+0]']
	-- 57 EOR [DP],Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH,AAL+YL->AAL']
	("000","011","10","000","00","01","00000101","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB','AAH+YH+AALCarry->AAH']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00110","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00110","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 58 CLI
	("010","000","00","100","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- ['[PBR:PC]->,ALU()->A', 'Flags', 'ALU()->X,Y', 'ALU()->A'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 59 EOR ABS,Y
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB'] 
	("001","000","00","000","00","01","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00110","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00110","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 5A PHY
	("110","000","00","000","00","00","00000000","000","000","011","00","000000","00000","00","000","00"),-- []
	("000","010","00","000","00","00","00000000","000","011","011","00","010000","00000","10","101","10"),-- ['YH->[00:SP]', 'SP--']
	("010","010","00","000","00","00","00000000","000","011","011","00","010000","00000","01","101","10"),-- ['YL->[00:SP]', 'SP--']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 5B TCD
	("010","000","00","001","00","00","00000000","000","000","000","01","000010","00001","00","000","00"),-- ['ALU(A)->D', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 5C JMP LONG
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++'] 
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++'] 
	("010","000","00","000","00","00","00000000","110","000","000","10","000000","00000","00","000","01"),-- ['[PBR:PC]->PBR', 'AA->PC'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 5D EOR ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("001","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00110","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00110","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 5E LSR ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("110","101","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[AB:AA+0]->TL'] 
	("000","101","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[AB:AA+1]->TH'] 
	("110","101","01","001","10","00","00000000","000","000","000","00","000100","01011","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","101","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[AB:AA+1]']
	("010","101","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[AB:AA+0]']
	-- 5F EOR LONG,X
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","000","00","000","00","00","00000101","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'PC++', 'AAH+XH/YH+AALCarry->AAH']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00110","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00110","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 60 RTS
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- ['']
	("000","000","00","000","00","00","00000000","000","001","000","00","000000","00000","00","000","00"),-- ['SP++']
	("000","010","00","000","00","00","00000000","000","001","000","00","000000","00000","00","000","10"),-- ['[00:SP]->DR', 'SP++']
	("000","010","00","000","00","00","00000000","010","000","000","00","000000","00000","00","000","10"),-- ['[00:SP]:DR->PC']
	("010","010","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","00"),-- ['PC++']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 61 ADC (DP,X)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00111","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']  
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00111","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 62 PER
	("000","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->TL', 'PC++'] 
	("000","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->TH', 'PC++'] 
	("000","000","00","000","00","00","01101100","000","000","000","00","000000","00000","00","000","00"),-- ['PC+Offset->AA'] 
	("000","010","00","000","00","00","00000000","000","011","000","00","000000","00000","10","011","10"),-- ['AAH->[00:SP]', 'SP--'] 
	("010","010","00","000","00","00","00000000","000","011","000","00","000000","00000","01","011","10"),-- ['AAL->[00:SP]', 'SP--'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 63 ADC S
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00111","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00111","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 64 STZ DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","000","00","00","00000000","000","000","000","00","000000","00000","01","111","10"),-- ['0->[00:DX+0]']
	("010","011","01","000","00","00","00000000","000","000","000","00","000000","00000","10","111","10"),-- ['0->[00:DX+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 65 ADC DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00111","01","000","10"),-- ['[00:DX+0]->A']   
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00111","10","000","10"),-- ['[00:DX+1]->A'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 66 ROR DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("110","011","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:DX+0]->TL'] 
	("000","011","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[00:DX+1]->TH'] 
	("110","011","01","001","10","00","00000000","000","000","000","00","000100","01101","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","011","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[00:DX+1]']
	("010","011","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[00:DX+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 67 ADC [DP]
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("000","011","10","000","00","00","00000001","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00111","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00111","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 68 PLA
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- 
	("000","000","00","000","00","00","00000000","000","001","000","00","000000","00000","00","000","00"),-- ['SP++']
	("100","010","00","001","00","00","00000000","000","010","101","00","000000","00000","01","000","10"),-- ['ALU([00:SP])->REGL', 'SP++']
	("010","010","00","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([00:SP])->REGH', 'SP++']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 69 ADC IMM
	("100","000","00","001","00","00","00000000","001","000","101","00","000000","00111","01","000","01"),-- ['ALU([PBR:PC])->AL', '[PBR:PC]->DR', 'PC++', 'Flags'] 
	("010","000","00","001","00","00","00000000","001","000","101","00","000001","00111","10","000","01"),-- ['ALU([PBR:PC]:DR)->A', 'PC++', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 6A ROR A
	("010","000","00","001","00","00","00000000","000","000","101","00","000010","01101","11","000","00"),-- ['ALU(REG+1)->REG', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 6B RTL
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- ['']
	("000","000","00","000","00","00","00000000","000","001","000","00","000000","00000","00","000","00"),-- ['SP++']
	("000","010","00","000","00","00","00000000","000","001","000","00","000000","00000","00","000","10"),-- ['[00:SP]->DR', 'SP++']
	("000","010","00","000","00","00","00000000","010","001","000","00","000000","00000","00","000","10"),-- ['[00:SP]:DR->PC', 'SP++']
	("010","010","00","000","00","00","00000000","001","000","000","10","000000","00000","00","000","10"),-- ['[00:SP]->PBR', 'PC++']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 6C JMP (ABS)
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++'] 
	("000","110","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:AA+0]->DR'] 
	("010","110","01","000","00","00","00000000","010","000","000","00","000000","00000","00","000","10"),-- ['[00:AA+1]:DR->PC'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 6D ADC ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00111","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags'] 
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00111","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 6E ROR ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++'] 
	("110","001","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[DBR:AA+0]->TL'] 
	("000","001","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[DBR:AA+1]->TH'] 
	("110","001","01","001","10","00","00000000","000","000","000","00","000100","01101","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","001","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[DBR:AA+1]']
	("010","001","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[DBR:AA+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 6F ADC LONG
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("000","000","00","000","00","00","00000001","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'PC++']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00111","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00111","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 70 BVS
	("010","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->DR', 'PC++'] 
	("011","000","00","000","00","00","00000000","100","000","000","00","000000","00000","00","000","00"),-- ['PC+DR->PC']
	("010","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- [] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 71 ADC (DP),Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB']
	("001","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL ']
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00111","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00111","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 72 ADC (DP)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- [00:DX+0]->AAL
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- [00:DX+1]->AAH
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00111","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']  
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00111","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 73 ADC (S),Y
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB'] 
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL']
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00111","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00111","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 74 STZ DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("100","011","00","000","00","00","00000000","000","000","000","00","000000","00000","01","111","10"),-- ['0->[00:DX+0]']
	("010","011","01","000","00","00","00000000","000","000","000","00","000000","00000","10","111","10"),-- ['0->[00:DX+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 75 ADC DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+Carry->DX'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00111","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00111","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 76 ROR DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("110","011","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:DX+0]->TL'] 
	("000","011","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[00:DX+1]->TH'] 
	("110","011","01","001","10","00","00000000","000","000","000","00","000100","01101","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","011","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[00:DX+1]']
	("010","011","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[00:DX+0]']
	-- 77 ADC [DP],Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL']
	("000","011","10","000","00","01","00000101","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB', 'AAH+YH+AALCarry->AAH']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00111","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00111","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 78 SEI
	("010","000","00","100","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- ['[PBR:PC]->,ALU()->A', 'Flags', 'ALU()->X,Y', 'ALU()->A'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 79 ADC ABS,Y
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("001","000","00","000","00","01","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00111","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00111","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 7A PLY
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("000","000","00","000","00","00","00000000","000","001","000","00","000000","00000","00","000","00"),-- ['SP++']
	("100","010","00","001","00","00","00000000","000","010","111","00","000000","00000","01","000","10"),-- ['ALU([00:SP])->YL', 'SP++']
	("010","010","00","001","00","00","00000000","000","000","111","00","000001","00001","10","000","10"),-- ['ALU([00:SP])->YH']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 7B TDC
	("010","000","00","001","00","00","00000000","000","000","101","00","011010","00001","11","000","00"),-- ['ALU(D)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 7C JMP (ABS,X)
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","000","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+Carry->AAH'] 
	("000","111","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","01"),-- ['[PBR:AA+0]->DR'] 
	("010","111","01","000","00","00","00000000","010","000","000","00","000000","00000","00","000","01"),-- ['[PBR:AA+1]:DR->PC'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 7D ADC ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("001","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH''] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00111","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00111","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 7E ROR ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("110","101","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[AB:AA+0]->TL'] 
	("000","101","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[AB:AA+1]->TH'] 
	("110","101","01","001","10","00","00000000","000","000","000","00","000100","01101","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","101","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[AB:AA+1]']
	("010","101","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[AB:AA+0]']
	-- 7F ADC LONG,X
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL']  
	("000","000","00","000","00","00","00000101","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'PC++', 'AAH+XH/YH+AALCarry->AAH']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00111","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00111","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 80 BRA
	("000","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->DL', 'PC++'] 
	("011","000","00","000","00","00","00000000","100","000","000","00","000000","00000","00","000","00"),-- ['PC+DL->PC']
	("010","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- [] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 81 STA (DP,X)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("100","001","00","000","00","00","00000000","000","000","000","00","000010","00000","01","101","10"),-- ['A->[DBR:AA+0]']
	("010","001","01","000","00","00","00000000","000","000","000","00","000010","00000","10","101","10"),-- ['B->[DBR:AA+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 82 BRL
	("000","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","01101100","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]:DL->AA', 'PC++'] 
	("010","000","00","000","00","00","00000000","011","000","000","00","000000","00000","00","000","00"),-- ['PC+Offset->PC'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 83 STA S
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['SPH+Carry->DH']
	("100","011","00","000","00","00","00000000","000","000","001","00","000010","00000","01","101","10"),-- ['REGL->[00:DX+0]']
	("010","011","01","000","00","00","00000000","000","000","001","00","000010","00000","10","101","10"),-- ['REGH->[00:DX+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 84 STY DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","000","00","00","00000000","000","000","011","00","010010","00000","01","101","10"),-- REGL->[00:DX+0]
	("010","011","01","000","00","00","00000000","000","000","011","00","010010","00000","10","101","10"),-- REGH->[00:DX+1]
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 85 STA DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","000","00","00","00000000","000","000","001","00","000010","00000","01","101","10"),-- REGL->[00:DX+0]
	("010","011","01","000","00","00","00000000","000","000","001","00","000010","00000","10","101","10"),-- REGH->[D00:X+1]
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 86 STX DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","000","00","00","00000000","000","000","010","00","001010","00000","01","101","10"),-- REGL->[00:DX+0]
	("010","011","01","000","00","00","00000000","000","000","010","00","001010","00000","10","101","10"),-- REGH->[00:DX+1]
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 87 STA [DP]
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("000","011","10","000","00","00","00000001","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB']
	("100","101","00","000","00","00","00000000","000","000","001","00","000010","00000","01","101","10"),-- ['REGL->[AB:AA+0]']
	("010","101","01","000","00","00","00000000","000","000","001","00","000010","00000","10","101","10"),-- ['REGH->[AB:AA+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 88 DEY
	("010","000","00","001","00","00","00000000","000","000","111","00","010010","00010","11","000","00"),-- ['ALU(Y)->Y', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 89 BIT IMM
	("100","000","00","111","00","00","00000000","001","000","001","00","000000","01001","01","000","01"),-- ['ALU([PBR:PC])', '[PBR:PC]->DR', 'PC++', 'Flags']   
	("010","000","00","111","00","00","00000000","001","000","001","00","000001","01001","10","000","01"),-- ['ALU([PBR:PC]:DR)', 'PC++', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 8A TXA
	("010","000","00","001","00","00","00000000","000","000","101","00","001010","00000","11","000","00"),-- ['ALU(X)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 8B PHB
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("010","010","00","000","00","00","00000000","000","011","000","00","111010","00000","01","101","10"),-- ['DBR->[00:SP]', 'SP--']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 8C STY ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","000","00","00","00000000","000","000","011","00","010010","00000","01","101","10"),-- ['REGL->[DBR:AA+0]']
	("010","001","01","000","00","00","00000000","000","000","011","00","010010","00000","10","101","10"),-- ['REGH->[DBR:AA+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 8D STA ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","000","00","00","00000000","000","000","001","00","000010","00000","01","101","10"),-- ['REGL->[DBR:AA+0]']
	("010","001","01","000","00","00","00000000","000","000","001","00","000010","00000","10","101","10"),-- ['REGH->[DBR:AA+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 8E STX ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++'] 
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","000","00","00","00000000","000","000","010","00","001010","00000","01","101","10"),-- ['REGL->[DBR:AA+0]']
	("010","001","01","000","00","00","00000000","000","000","010","00","001010","00000","10","101","10"),-- ['REGH->[DBR:AA+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 8F STA LONG
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("000","000","00","000","00","00","00000001","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'PC++']
	("100","101","00","000","00","00","00000000","000","000","001","00","000010","00000","01","101","10"),-- ['REGL->[AB:AA+0]']
	("010","101","01","000","00","00","00000000","000","000","001","00","000010","00000","10","101","10"),-- ['REGH->[AB:AA+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 90 BCC
	("010","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->DR', 'PC++'] 
	("011","000","00","000","00","00","00000000","100","000","000","00","000000","00000","00","000","00"),-- ['PC+DR->PC']
	("010","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- [] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 91 STA (DP),Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB']
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL ']
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","000","00","00","00000000","000","000","001","00","000010","00000","01","101","10"),-- ['A->[AB:AA+0]']
	("010","101","01","000","00","00","00000000","000","000","001","00","000010","00000","10","101","10"),-- ['B->[AB:AA+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 92 STA (DP)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("100","001","00","000","00","00","00000000","000","000","001","00","000010","00100","01","101","10"),-- ['A->[DBR:AA+0]']
	("010","001","01","000","00","00","00000000","000","000","001","00","000010","00000","10","101","10"),-- ['B->[DBR:AA+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 93 STA (S),Y
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['SPH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB'] 
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL']
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","000","00","00","00000000","000","000","001","00","000010","00000","01","101","10"),-- ['REGL->[AB:AA+0]']
	("010","101","01","000","00","00","00000000","000","000","001","00","000010","00000","10","101","10"),-- ['REGH->[AB:AA+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 94 STY DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("100","011","00","000","00","00","00000000","000","000","011","00","010010","00000","01","101","10"),-- ['REGL->[00:DX+0]']
	("010","011","01","000","00","00","00000000","000","000","011","00","010010","00000","10","101","10"),-- ['REGH->[00:DX+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 95 STA DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("100","011","00","000","00","00","00000000","000","000","001","00","000010","00000","01","101","10"),-- ['REGL->[00:DX+0]']
	("010","011","01","000","00","00","00000000","000","000","001","00","000010","00000","10","101","10"),-- ['REGH->[00:DX+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 96 STX DP,Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","000","00","000","00","01","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+Y->DX']
	("100","011","00","000","00","00","00000000","000","000","010","00","001010","00000","01","101","10"),-- ['REGL->[00:DX+0]']
	("010","011","01","000","00","00","00000000","000","000","010","00","001010","00000","10","101","10"),-- ['REGH->[00:DX+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 97 STA [DP],Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH,AAL+YL->AAL']
	("000","011","10","000","00","01","00000101","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB','AAH+YH+AALCarry->AAH']
	("100","101","00","000","00","00","00000000","000","000","001","00","000010","00000","01","101","10"),-- ['REGL->[AB:AA+0]']
	("010","101","01","000","00","00","00000000","000","000","001","00","000010","00000","10","101","10"),-- ['REGH->[AB:AA+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 98 TYA
	("010","000","00","001","00","00","00000000","000","000","101","00","010010","00000","11","000","00"),-- ['ALU(Y)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 99 STA ABS,Y
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB'] 
	("000","000","00","000","00","01","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","000","00","00","00000000","000","000","001","00","000010","00000","01","101","10"),-- ['A->[AB:AA+0]'] 
	("010","101","01","000","00","00","00000000","000","000","001","00","000010","00000","10","101","10"),-- ['B->[AB:AA+1]'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 9A TXS
	("010","000","00","000","00","00","00000000","000","101","000","00","000000","00000","00","000","00"),-- ['X->S'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 9B TXY
	("010","000","00","001","00","00","00000000","000","000","111","00","001010","00000","11","000","00"),-- ['ALU(X)->Y', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 9C STZ ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","000","00","00","00000000","000","000","000","00","000000","00000","01","111","10"),-- ALU(0)->[DBR:AA+0]
	("010","001","01","000","00","00","00000000","000","000","000","00","000000","00000","10","111","10"),-- ALU(0)->[DBR:AA+1]
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 9D STA ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","000","00","00","00000000","000","000","001","00","000010","00000","01","101","10"),-- ['A->[AB:AA+0]']
	("010","101","01","000","00","00","00000000","000","000","001","00","000010","00000","10","101","10"),-- ['B->[AB:AA+1]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 9E STZ ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","000","00","00","00000000","000","000","000","00","000000","00000","01","111","10"),-- ALU(0)->[AB:AA+0]
	("010","101","01","000","00","00","00000000","000","000","000","00","000000","00000","10","111","10"),-- ALU(0)->[AB:AA+1]
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- 9F STA LONG,X
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","000","00","000","00","00","00000101","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'PC++', 'AAH+XH/YH+AALCarry->AAH']
	("100","101","00","000","00","00","00000000","000","000","001","00","000010","00000","01","101","10"),-- ['A->[AB:AA+0]'] 
	("010","101","01","000","00","00","00000000","000","000","001","00","000010","00000","10","101","10"),-- ['B->[AB:AA+1]'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	--A0 LDY IMM
	("100","000","00","001","00","00","00000000","001","000","111","00","000000","00000","01","000","01"),-- ['ALU([PBR:PC])->YL', '[PBR:PC]->DR', 'PC++', 'Flags'] 
	("010","000","00","001","00","00","00000000","001","000","111","00","000001","00001","10","000","01"),-- ['ALU([PBR:PC]:DR)->Y', 'PC++', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- A1 LDA (DP,X)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00000","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']  
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- A2 LDX IMM
	("100","000","00","001","00","00","00000000","001","000","110","00","000000","00000","01","000","01"),-- ['ALU([PBR:PC])->XL', '[PBR:PC]->DR', 'PC++', 'Flags']  
	("010","000","00","001","00","00","00000000","001","000","110","00","000001","00001","10","000","01"),-- ['ALU([PBR:PC]:DR)->X', 'PC++', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- A3 LDA S
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00000","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']   
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- A4 LDY DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("100","011","00","001","00","00","00000000","000","000","111","00","000000","00000","01","000","10"),-- ['ALU([00:DX+0]->YL', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","111","00","000001","00001","10","000","10"),-- ['ALU([00:DX+1]->Y', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- A5 LDA DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00000","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']   
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- A6 LDX DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","110","00","000000","00000","01","000","10"),-- ['ALU([00:DX+0]->XL', '[00:DX+0]->DR', 'Flags'] 
	("010","011","01","001","00","00","00000000","000","000","110","00","000001","00001","10","000","10"),-- ['ALU([00:DX+1]->X', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- A7 LDA [DP]
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("000","011","10","000","00","00","00000001","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']   
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- A8 TAY
	("010","000","00","001","00","00","00000000","000","000","111","00","000010","00000","11","000","00"),-- ['ALU(A)->Y', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- A9 LDA IMM
	("100","000","00","001","00","00","00000000","001","000","101","00","000000","00000","01","000","01"),-- ['ALU([PBR:PC])->AL', '[PBR:PC]->DR', 'PC++', 'Flags'] 
	("010","000","00","001","00","00","00000000","001","000","101","00","000001","00001","10","000","01"),-- ['ALU([PBR:PC]:DR)->A', 'PC++', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- AA TAX
	("010","000","00","001","00","00","00000000","000","000","110","00","000010","00000","11","000","00"),-- ['ALU(A)->X', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- AB PLB
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("000","000","00","000","00","00","00000000","000","001","000","00","000000","00000","00","000","00"),-- ['SP++']
	("010","010","00","001","00","00","00000000","000","000","000","11","000000","00000","00","000","10"),-- ['ALU([00:SP])->DBR']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- AC LDY ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","001","00","00","00000000","000","000","111","00","000000","00000","01","000","10"),-- ['ALU([DBR:AA+0])->YL', '[DBR:AA+0]->DR', 'Flags']
	("010","001","01","001","00","00","00000000","000","000","111","00","000001","00001","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->Y', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- AD LDA ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00000","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- AE LDX ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","001","00","00","00000000","000","000","110","00","000000","00000","01","000","10"),-- ['ALU([DBR:AA+0])->XL', '[DBR:AA+0]->DR', 'Flags']
	("010","001","01","001","00","00","00000000","000","000","110","00","000001","00001","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->X', 'Flags']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- AF LDA LONG
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("000","000","00","000","00","00","00000001","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'PC++']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- B0 BCS
	("010","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->DR', 'PC++'] 
	("011","000","00","000","00","00","00000000","100","000","000","00","000000","00000","00","000","00"),-- ['PC+DR->PC']
	("010","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- [] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- B1 LDA (DP),Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB']
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL ']
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- B2 LDA (DP)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH ']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","00000","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags'] 
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- B3 LDA (S),Y
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['SPH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB'] 
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL'] 
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']   
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- B4 LDY DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- [DX+X->DX]
	("100","011","00","001","00","00","00000000","000","000","111","00","000000","00000","01","000","10"),-- ['ALU([00:DX+0]->YL', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","111","00","000001","00001","10","000","10"),-- ['ALU([00:DX+1]->Y', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- B5 LDA DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+Carry->DX'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","00000","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- B6 LDX DP,Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+Carry->DX'] 
	("000","000","00","000","00","01","10010000","000","000","000","00","000000","00000","00","000","00"),-- [DX+Y->DX]
	("100","011","00","001","00","00","00000000","000","000","110","00","000000","00000","01","000","10"),-- ['ALU([00:DX+0]->XL', '[00:DX+0]->DR', 'Flags'] 
	("010","011","01","001","00","00","00000000","000","000","110","00","000001","00001","10","000","10"),-- ['ALU([00:DX+1]->X', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- B7 LDA [DP],Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH,AAL+YL->AAL']
	("000","011","10","000","00","01","00000101","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB','AAH+YH+AALCarry->AAH']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']   
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- B8 CLV
	("010","000","00","100","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- ['[PC]->,ALU()->A', 'Flags', 'ALU()->X,Y', 'ALU()->A'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- B9 LDA ABS,Y
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("001","000","00","000","00","01","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- BA TSX
	("010","000","00","001","00","00","00000000","000","000","110","00","101010","00001","11","000","00"),-- ['ALU(SP)->X', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- BB TYX
	("010","000","00","001","00","00","00000000","000","000","110","00","010010","00000","11","000","00"),-- ['ALU(Y)->X', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- BC LDY ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("001","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","111","00","000000","00000","01","000","10"),-- ['ALU([AB:AA+0])->YL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","111","00","000001","00001","10","000","10"),-- ['ALU([AB:AA+1])->Y', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- BD LDA ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("001","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- BE LDX ABS,Y
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("001","000","00","000","00","01","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL']  
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","110","00","000000","00000","01","000","10"),-- ['ALU([AB:AA+0])->XL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","110","00","000001","00001","10","000","10"),-- ['ALU([AB:AA+1])->X', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- BF LDA LONG,X
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","000","00","000","00","00","00000101","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'PC++', 'AAH+XH/YH+AALCarry->AAH']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","00000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","00001","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- C0 CPY IMM
	("100","000","00","001","00","00","00000000","001","000","011","00","010000","10000","01","000","01"),-- ['ALU([PBR:PC])', '[PBR:PC]->DR', 'PC++', 'Flags'] 
	("010","000","00","001","00","00","00000000","001","000","011","00","010001","10000","10","000","01"),-- ['ALU([PBR:PC]:DR)', 'PC++', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- C1 CMP (DP,X)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("100","001","00","001","00","00","00000000","000","000","001","00","000000","10000","01","000","10"),-- ['ALU([AB:AA+0])', '[AB:AA+0]->DR', 'Flags']   
	("010","001","01","001","00","00","00000000","000","000","001","00","000001","10000","10","000","10"),-- ['ALU([AB:AA+1])', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- C2 REP
	("000","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- [[PBR:PC]->DR', 'PC++'] 
	("010","000","00","110","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- ['Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- C3 CMP S
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['SPH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","001","00","000000","10000","01","000","10"),-- ['ALU([00:DX+0]', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","001","00","000001","10000","10","000","10"),-- ['ALU([00:DX+1]', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- C4 CPY DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","011","00","010000","10000","01","000","10"),-- ['ALU([00:DX+0]', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","011","00","010001","10000","10","000","10"),-- ['ALU([00:DX+1]', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- C5 CMP DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","001","00","000000","10000","01","000","10"),-- ['ALU([00:DX+0]', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","001","00","000001","10000","10","000","10"),-- ['ALU([00:DX+1]', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- C6 DEC DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("110","011","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:DX+0]->TL'] 
	("000","011","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[00:DX+1]->TH'] 
	("110","011","01","001","10","00","00000000","000","000","000","00","100010","00010","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","011","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[00:DX+1]']
	("010","011","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[00:DX+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- C7 CMP [DP]
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("000","011","10","000","00","00","00000001","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB']
	("100","101","00","001","00","00","00000000","000","000","001","00","000000","10000","01","000","10"),-- ['ALU([AB:AA+0])', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","001","00","000001","10000","10","000","10"),-- ['ALU([AB:AA+1])', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- C8 INY
	("010","000","00","001","00","00","00000000","000","000","111","00","010010","00011","11","000","00"),-- ['ALU(Y+1)->Y', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- C9 CMP IMM
	("100","000","00","001","00","00","00000000","001","000","001","00","000000","10000","01","000","01"),-- ['ALU([PBR:PC])', '[PBR:PC]->DR', 'PC++', 'Flags'] 
	("010","000","00","001","00","00","00000000","001","000","001","00","000001","10000","10","000","01"),-- ['ALU([PBR:PC]:DR)', 'PC++', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- CA DEX
	("010","000","00","001","00","00","00000000","000","000","110","00","001010","00010","11","000","00"),-- ['ALU(X-1)->X', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- CB WAI
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("010","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- CC CPY ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","001","00","00","00000000","000","000","011","00","010000","10000","01","000","10"),-- ['ALU([DBR:AA+0])', '[DBR:AA+0]->DR', 'Flags']
	("010","001","01","001","00","00","00000000","000","000","011","00","010001","10000","10","000","10"),-- ['ALU([DBR:AA+1]:DR)', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- CD CMP ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","001","00","00","00000000","000","000","001","00","000000","10000","01","000","10"),-- ['ALU([DBR:AA+0])', '[DBR:AA+0]->DR', 'Flags']
	("010","001","01","001","00","00","00000000","000","000","001","00","000001","10000","10","000","10"),-- ['ALU([DBR:AA+1]:DR)', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- CE DEC ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++'] 
	("110","001","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[DBR:AA+0]->TL'] 
	("000","001","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[DBR:AA+1]->TH'] 
	("110","001","01","001","10","00","00000000","000","000","000","00","100010","00010","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","001","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[DBR:AA+1]']
	("010","001","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[DBR:AA+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- CF CMP LONG
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("000","000","00","000","00","00","00000001","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'PC++']
	("100","101","00","001","00","00","00000000","000","000","001","00","000000","10000","01","000","10"),-- ['ALU([AB:AA+0])', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","001","00","000001","10000","10","000","10"),-- ['ALU([AB:AA+1])', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- D0 BNE
	("010","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->DR', 'PC++'] 
	("011","000","00","000","00","00","00000000","100","000","000","00","000000","00000","00","000","00"),-- ['PC+DR->PC']
	("010","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- [] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- D1 CMP (DP),Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB']
	("001","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL ']
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","001","00","000000","10000","01","000","10"),-- ['ALU([AB:AA+0])', '[AB:AA+0]->DR', 'Flags']   
	("010","101","01","001","00","00","00000000","000","000","001","00","000001","10000","10","000","10"),-- ['ALU([AB:AA+1])', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- D2 CMP (DP)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("100","001","00","001","00","00","00000000","000","000","001","00","000000","10000","01","000","10"),-- ['ALU([DBR:AA+0])', '[DBR:AA+0]->DR', 'Flags']
	("010","001","01","001","00","00","00000000","000","000","001","00","000001","10000","10","000","10"),-- ['ALU([DBR:AA+1]:DR)', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- D3 CMP (S),Y
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['SPH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR+AAHCarry->AB']
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL']
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","001","00","000000","10000","01","000","10"),-- ['ALU([AB:AA+0])', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","001","00","000001","10000","10","000","10"),-- ['ALU([AB:AA+1])', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- D4 PEI
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("000","010","00","000","00","00","00000000","000","011","000","00","000000","00000","10","011","10"),-- ['AAH->[00:SP]', 'SP--'] 
	("010","010","00","000","00","00","00000000","000","011","000","00","000000","00000","01","011","10"),-- ['AAL->[00:SP]', 'SP--'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- D5 CMP DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+Carry->DX'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("100","011","00","001","00","00","00000000","000","000","001","00","000000","10000","01","000","10"),-- ['ALU([00:DX+0]', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","001","00","000001","10000","10","000","10"),-- ['ALU([00:DX+1]', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- D6 DEC DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("110","011","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:DX+0]->TL'] 
	("000","011","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[00:DX+1]->TH'] 
	("110","011","01","001","10","00","00000000","000","000","000","00","100010","00010","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","011","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[DX+1]']
	("010","011","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[DX+0]']
	-- D7 CMP [DP],Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH,AAL+YL->AAL']
	("000","011","10","000","00","01","00000101","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB','AAH+YH+AALCarry->AAH']
	("100","101","00","001","00","00","00000000","000","000","001","00","000000","10000","01","000","10"),-- ['ALU([AB:AA+0])', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","001","00","000001","10000","10","000","10"),-- ['ALU([AB:AA+1])', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- D8 CLD
	("010","000","00","100","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- ['[PC]->,ALU()->A', 'Flags', 'ALU()->X,Y', 'ALU()->A'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- D9 CMP ABS,Y
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("001","000","00","000","00","01","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","001","00","000000","10000","01","000","10"),-- ['ALU([AB:AA+0])', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","001","00","000001","10000","10","000","10"),-- ['ALU([AB:AA+1])', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- DA PHX
	("110","000","00","000","00","00","00000000","000","000","010","00","000000","00000","00","000","00"),-- []
	("000","010","00","000","00","00","00000000","000","011","010","00","001000","00000","10","101","10"),-- ['XH->[00:SP]', 'SP--']
	("010","010","00","000","00","00","00000000","000","011","010","00","001000","00000","01","101","10"),-- ['XL->[00:SP]', 'SP--']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- DB STP
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("010","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- DC JMP [ABS]
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++'] 
	("000","110","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:AA+0]->DL']
	("000","110","01","000","00","00","00000000","010","000","000","00","000000","00000","00","000","10"),-- ['[00:AA+1]:DL->PC'] 
	("010","110","10","000","00","00","00000000","000","000","000","10","000000","00000","00","000","10"),-- ['[00:AA+2]->PBR'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- DD CMP ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("001","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","001","00","000000","10000","01","000","10"),-- ['ALU([AB:AA+0])', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","001","00","000001","10000","10","000","10"),-- ['ALU([AB:AA+1])', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- DE DEC ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("110","101","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[AB:AA+0]->TL'] 
	("000","101","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[AB:AA+1]->TH'] 
	("110","101","01","001","10","00","00000000","000","000","000","00","100010","00010","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","101","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[AB:AA+1]']
	("010","101","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[AB:AA+0]']
	-- DF CMP LONG,X
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","000","00","000","00","00","00000101","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'PC++', 'AAH+XH/YH+AALCarry->AAH']
	("100","101","00","001","00","00","00000000","000","000","001","00","000000","10000","01","000","10"),-- ['ALU([AB:AA+0])', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","001","00","000001","10000","10","000","10"),-- ['ALU([AB:AA+1])', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- E0 CPX IMM
	("100","000","00","001","00","00","00000000","001","000","010","00","001000","10000","01","000","01"),-- ['ALU([PBR:PC])', '[PBR:PC]->DR', 'PC++', 'Flags'] 
	("010","000","00","001","00","00","00000000","001","000","010","00","001001","10000","10","000","01"),-- ['ALU([PBR:PC]:DR)', 'PC++', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- E1 SBC (DP,X)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","01000","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","01000","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- E2 SEP
	("000","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]-DR', 'PC++'] 
	("010","000","00","110","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- ['Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- E3 SBC S
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['SPH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","01000","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","01000","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- E4 CPX DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","010","00","001000","10000","01","000","10"),-- ['ALU([00:DX+0]', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","010","00","001001","10000","10","000","10"),-- ['ALU([00:DX+1]', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- E5 SBC DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","01000","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","01000","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- E6 INC DP
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("110","011","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:DX+0]->TL'] 
	("000","011","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[00:DX+1]->TH'] 
	("110","011","01","001","10","00","00000000","000","000","000","00","100010","00011","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","011","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[00:DX+1]']
	("010","011","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[00:DX+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- E7 SBC [DP]
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("000","011","10","000","00","00","00000001","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","01000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","01000","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- E8 INX
	("010","000","00","001","00","00","00000000","000","000","110","00","001010","00011","11","000","00"),-- ['ALU(REG+1)->REG', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- E9 SBC IMM
	("100","000","00","001","00","00","00000000","001","000","101","00","000000","01000","01","000","01"),-- ['ALU([PBR:PC])->AL', '[PBR:PC]->DR', 'PC++', 'Flags']   
	("010","000","00","001","00","00","00000000","001","000","101","00","000001","01000","10","000","01"),-- ['ALU([PBR:PC]:DR)->A', 'PC++', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- EA NOP
	("010","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- []
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- EB XBA
	("000","000","00","000","00","00","00000000","000","000","101","00","000000","00000","11","000","00"),-- ['B:A->C']
	("010","000","00","001","00","00","00000000","000","000","001","00","000010","00000","01","000","00"),-- ['Flags']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- EC CPX ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","001","00","00","00000000","000","000","010","00","001000","10000","01","000","10"),-- ['ALU([DBR:AA+0])', '[DBR:AA+0]->DR', 'Flags']
	("010","001","01","001","00","00","00000000","000","000","010","00","001001","10000","10","000","10"),-- ['ALU([DBR:AA+1]:DR)', 'Flags']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- ED SBC ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","01000","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","01000","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- EE INC ABS
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++'] 
	("110","001","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[DBR:AA+0]->TL'] 
	("000","001","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[DBR:AA+1]->TH'] 
	("110","001","01","001","10","00","00000000","000","000","000","00","100010","00011","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","001","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[DBR:AA+1]']
	("010","001","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[DBR:AA+0]']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- EF SBC LONG
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("000","000","00","000","00","00","00000001","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'PC++']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","01000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","01000","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- F0 BEQ
	("010","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->DR', 'PC++'] 
	("011","000","00","000","00","00","00000000","100","000","000","00","000000","00000","00","000","00"),-- ['PC+DR->PC']
	("010","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- [] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- F1 SBC (DP),Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB']
	("001","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL ']
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","01000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","01000","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- F2 SBC (DP)
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH'] 
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","00","00001000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH']
	("100","001","00","001","00","00","00000000","000","000","101","00","000000","01000","01","000","10"),-- ['ALU([DBR:AA+0])->AL', '[DBR:AA+0]->DR', 'Flags']
	("010","001","01","001","00","00","00000000","000","000","101","00","000001","01000","10","000","10"),-- ['ALU([DBR:AA+1]:DR)->A', 'Flags']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- F3 SBC (S),Y
	("000","000","00","000","00","00","10110111","001","000","000","00","000000","00000","00","000","01"),-- ['SPL+[PBR:PC]->DL', 'PC++'] 
	("000","000","00","000","00","00","00011011","000","000","000","00","000000","00000","00","000","00"),-- ['SPH+Carry->DH'] 
	("000","011","00","000","00","00","01000011","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL', 'DBR->AB'] 
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH', 'AAL+YL->AAL'] 
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","01000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","01000","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- F4 PEA
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00001000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++']
	("000","010","00","000","00","00","00000000","000","011","000","00","000000","00000","10","011","10"),-- ['AAH->[00:SP]', 'SP--'] 
	("010","010","00","000","00","00","00000000","000","011","000","00","000000","00000","01","011","10"),-- ['AAL->[00:SP]', 'SP--'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- F5 SBC DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+Carry->DX'] 
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("100","011","00","001","00","00","00000000","000","000","101","00","000000","01000","01","000","10"),-- ['ALU([00:DX+0])->AL', '[00:DX+0]->DR', 'Flags']  
	("010","011","01","001","00","00","00000000","000","000","101","00","000001","01000","10","000","10"),-- ['ALU([00:DX+1]:DR)->A', 'Flags'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- F6 INC DP,X
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","000","00","000","00","00","10010000","000","000","000","00","000000","00000","00","000","00"),-- ['DX+X->DX']
	("110","011","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[00:DX+0]->TL'] 
	("000","011","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[00:DX+1]->TH'] 
	("110","011","01","001","10","00","00000000","000","000","000","00","100010","00011","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","011","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[00:DX+1]']
	("010","011","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[00:DX+0]']
	-- F7 SBC [DP],Y
	("101","000","00","000","00","00","10110100","001","000","000","00","000000","00000","00","000","01"),-- ['DL+[PBR:PC]->DL', 'PC++']
	("000","000","00","000","00","00","00011000","000","000","000","00","000000","00000","00","000","00"),-- ['DH+Carry->DH']
	("000","011","00","000","00","00","01000000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+0]->AAL']
	("000","011","01","000","00","01","00101000","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+1]->AAH,AAL+YL->AAL']
	("000","011","10","000","00","01","00000101","000","000","000","00","000000","00000","00","000","10"),-- ['[00:DX+2]->AB','AAH+YH+AALCarry->AAH']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","01000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","01000","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- F8 SED
	("010","000","00","100","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- ['[PC]->,ALU()->A', 'Flags', 'ALU()->X,Y', 'ALU()->A'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- F9 SBC ABS,Y
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("001","000","00","000","00","01","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","01","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","01000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","01000","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- FA PLX
	("000","000","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- 
	("000","000","00","000","00","00","00000000","000","001","000","00","000000","00000","00","000","00"),-- ['SP++']
	("100","010","00","001","00","00","00000000","000","010","110","00","000000","00000","01","000","10"),-- ['ALU([00:SP])->REGL', 'SP++']
	("010","010","00","001","00","00","00000000","000","000","110","00","000001","00001","10","000","10"),-- ['ALU([00:SP])->REGH']
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- FB XCE
	("010","000","00","101","00","00","00000000","000","000","000","00","000000","00000","00","000","00"),-- ['[PC]->,ALU()->A', 'Flags', 'ALU()->X,Y', 'ALU()->A'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- FC JSR (ABS,X)
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","010","00","000","00","00","00000000","000","011","000","00","000000","00000","10","010","10"),-- ['PCH->[00:SP]', 'SP--'] 
	("000","010","00","000","00","00","00000000","000","011","000","00","000000","00000","01","010","10"),-- ['PCL->[00:SP]', 'SP--'] 
	("000","000","00","000","00","00","00101000","000","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'AAL+XL/YL->AAL'] 
	("000","000","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+Carry->AAH'] 
	("000","111","00","000","00","00","00000000","000","000","000","00","000000","00000","00","000","01"),-- ['[PBR:AA+0]->DR'] 
	("010","111","01","000","00","00","00000000","010","000","000","00","000000","00000","00","000","01"),-- ['[PBR:AA+1]:DR->PC'] 
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- FD SBC ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("001","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH']  
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","01000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","01000","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	-- FE INC ABS,X
	("000","000","00","000","00","00","01000011","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++', 'DBR->AB']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","101","00","000","00","00","00000100","000","000","000","00","000000","00000","00","000","00"),-- ['AAH+XH/YH+AALCarry->AAH'] 
	("110","101","00","000","01","00","00000000","000","000","000","00","000000","00000","01","000","10"),-- ['[AB:AA+0]->TL'] 
	("000","101","01","000","01","00","00000000","000","000","000","00","000000","00000","10","000","10"),-- ['[AB:AA+1]->TH'] 
	("110","101","01","001","10","00","00000000","000","000","000","00","100010","00011","11","000","00"),-- ['ALU(T)->T', 'Flags']
	("000","101","01","000","00","00","00000000","000","000","000","00","100000","00000","10","101","10"),-- ['TH->[AB:AA+1]']
	("010","101","00","000","00","00","00000000","000","000","000","00","100000","00000","01","101","10"),-- ['TL->[AB:AA+0]']
	-- FF SBC LONG,X
	("000","000","00","000","00","00","01000000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAL', 'PC++']
	("000","000","00","000","00","00","00101000","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AAH', 'PC++', 'AAL+XL/YL->AAL'] 
	("000","000","00","000","00","00","00000101","001","000","000","00","000000","00000","00","000","01"),-- ['[PBR:PC]->AB', 'PC++', 'AAH+XH/YH+AALCarry->AAH']
	("100","101","00","001","00","00","00000000","000","000","101","00","000000","01000","01","000","10"),-- ['ALU([AB:AA+0])->AL', '[AB:AA+0]->DR', 'Flags']  
	("010","101","01","001","00","00","00000000","000","000","101","00","000001","01000","10","000","10"),-- ['ALU([AB:AA+1]:DR)->A', 'Flags']  
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX"),
	("XXX","XXX","XX","XXX","XX","XX","XXXXXXXX","XXX","XXX","XXX","XX","XXXXXX","XXXXX","XX","XXX","XX")
	);
	

	type ALUCtrl_t is array(0 to 16) of ALUCtrl_r;
	constant ALU_TAB: ALUCtrl_t := (
	("100","100",'0','0'),-- 00000 LOAD 8BIT
	("100","100",'0','1'),-- 00001 LOAD 16BIT
	("110","100",'0','0'),-- 00010 DEC 
	("111","100",'0','0'),-- 00011 INC
	("100","000",'0','0'),-- 00100 ORA
	("100","001",'0','0'),-- 00101 AND
	("100","010",'0','0'),-- 00110 EOR
	("100","011",'0','0'),-- 00111 ADC
	("100","111",'1','0'),-- 01000 SBC
	("100","001",'1','0'),-- 01001 BIT
	("000","100",'0','0'),-- 01010 ASL
	("010","100",'0','0'),-- 01011 LSR
	("001","100",'0','0'),-- 01100 ROL
	("011","100",'0','0'),-- 01101 ROR
	("100","101",'0','0'),-- 01110 TRB
	("100","101",'1','0'),-- 01111 TSB
	("100","110",'0','0') -- 10000 CMP
	);
	
	signal MI    	: MicroInst_r;
	signal ALUFlags: ALUCtrl_r;

begin

	ALUFlags <= ALU_TAB(to_integer(unsigned(MI.ALUCtrl)));

	process(CLK, RST_N)
		variable STATE2 : unsigned(3 downto 0);
	begin
		if RST_N = '0' then
			MI <= ("000","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","11");
		elsif falling_edge(CLK) then
			STATE2 := STATE - 1;
			if EN = '1' then
				if STATE = "0000" then
					MI <= ("000","000","00","000","00","00","00000000","001","000","000","00","000000","00000","00","000","11");
				else
					MI <= M_TAB(to_integer(unsigned(IR) & STATE2(2 downto 0)));
				end if;
			end if;
		end if;
	end process;
	
	M <= (ALUFlags, MI.stateCtrl, MI.addrBus, MI.addrInc, MI.muxCtrl, MI.addrCtrl, MI.loadPC, MI.loadSP, 
			MI.regAXY, MI.loadP, MI.loadT, MI.loadDKB, MI.busCtrl, MI.byteSel, MI.outBus, MI.va);
	 
end rtl;